library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity clk_gen_p2 is
  port (
    END_SIM : in  std_logic;
    CLK     : out std_logic;
    RST_n   : out std_logic);
end clk_gen_p2 ;

architecture beh of clk_gen_p2  is

  constant Ts : time := 1.85 ns;
  constant Tp : time := 2 ns;
  
  signal CLK_i : std_logic;
  
begin  -- beh

  process
  begin  -- process
    if (CLK_i = 'U') then
      CLK_i <= '0';
    else
      CLK_i <= not(CLK_i);
    end if;
    wait for Ts/2;
  end process;

  CLK <= CLK_i and not(END_SIM);

  process
  begin  -- process
    RST_n <= '1';
    wait for Tp;
    RST_n <= '0';
    wait for 2*Ts;
    RST_n <= '1';
    wait;
  end process;

end beh;
